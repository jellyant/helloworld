//-- Fichero setbit.v
module setbit(output A);
wire A;
    
assign A = 1;
    
endmodule
